`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:30:06 01/20/2016 
// Design Name: 
// Module Name:    CLACell 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module CLACell(
		input a,
		input b,
		input c,
		output g,
		output p, 
		output s
	);
	
	assign g = a & b;
	assign p = a + b;
	assign s = a ^ b ^ c;

endmodule
